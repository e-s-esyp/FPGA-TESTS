module schema(
	CLOCK_50,
	pin_name1
);


input wire	CLOCK_50;
output wire	pin_name1;


assign	pin_name1 = CLOCK_50;




endmodule
