module con3(
	input wire [2:0] in,
	output wire [2:0] out
);

assign out = in;

endmodule
